----------------------------------------------------------------------------------
-- Ԫ�����ƣ�IDָ�������
-- ��������������һ��16λTHCO MIPSָ���������ָ�����������źźͼĴ�����š�
-- ��Ϊ������ָ�������Ϊ����߼���·�������������ı仯���仯������Ҫʱ���źź͸�λ�źš�
-- �˿�������
-- 	Insn		�������ָ��
-- 	Reg1		��һ�Ĵ����ı��
-- 	Reg2		�ڶ��Ĵ����ı��
--		RegDst	д�صļĴ������
--		Imm		������
-- 	Op1Src	ALU��һ��������Դ�Ŀ����ź�
-- 	Op2Src	ALU�ڶ���������Դ�Ŀ����ź�
-- 	AluOp		ALU�������
--		TWr		д��T�Ĵ��������ź�
--		Jcond		��ת��������
--		MemRd		�ڴ��ȡ�����ź�
--		MemWr		�ڴ�д������ź�
--		RegWr		д�ؼĴ��������ź�
--		Inval		�Ƿ�ָ���쳣
--		Priv		��Ȩָ���쳣
--		Lf			���м�
--		Degrade	�������м�
--		Int		INTָ��
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ID is
    Port ( Lf : in  STD_LOGIC;
			  Insn : in  STD_LOGIC_VECTOR(19 downto 0);
           Reg1 : out  STD_LOGIC_VECTOR(3 downto 0);
           Reg2 : out  STD_LOGIC_VECTOR(3 downto 0);
           RegDst : out  STD_LOGIC_VECTOR(3 downto 0);
			  Imm : out  STD_LOGIC_VECTOR(15 downto 0);
			  Op1Src : out  STD_LOGIC;
			  Op2Src : out  STD_LOGIC;
			  AluOp : out  STD_LOGIC_VECTOR(3 downto 0);
			  TWr : out  STD_LOGIC;
			  Jcond : out  STD_LOGIC_VECTOR(2 downto 0);
			  MemRd : out  STD_LOGIC;
			  MemWr : out  STD_LOGIC;
			  RegWr : out  STD_LOGIC;
			  Inval : out  STD_LOGIC;
			  Priv : out  STD_LOGIC;
			  Int : out  STD_LOGIC;
			  Degrade : out  STD_LOGIC);
end ID;

architecture Behavioral of ID is

begin
	process(Insn,Lf)
	begin
		-- ����Ϊ�������źŵ�Ĭ��ֵ����NOPָ����ͬ��
		Reg1 <= "1111"; -- Reg1 <= ZERO
		Reg2 <= "1111"; -- Reg2 <= ZERO
		RegDst <= "1111"; -- RegDst <= R0
		Imm <= "0000000000000000";
		Op1Src <= '0'; -- Data1
		Op2Src <= '0'; -- Data2
		AluOp <= "0000"; -- Add
		TWr <= '0'; -- No
		Jcond <= "000"; -- No
		MemRd <= '0'; -- No
		MemWr <= '0'; -- No
		RegWr <= '0'; -- No
		Inval <= '0'; -- No
		Priv <= '0'; -- No
		Degrade <= '0'; -- No
		Int <= '0'; -- No
		
		case Insn(19) is
			when '1' => -- CPU�쳣���ⳤָ��
				case Insn(18 downto 16) is
					when "000" => -- LI_ER
						RegDst <= "1011"; -- RegDst <= ER
						Imm <= Insn(15 downto 0);
						Op2Src <= '1'; -- Imm
						RegWr <= '1'; -- Yes
					when "001" => -- SW_ER
						Reg1 <= "1000"; -- Reg1 <= SP
						Reg2 <= "1011"; -- RegDst <= ER
						Imm <= Insn(15 downto 0);
						Op2Src <= '1'; -- Imm
						MemWr <= '1'; -- Yes
					when others => -- �Ƿ�ָ��
				end case;
			when others => -- ��ͨ16λָ��
				case Insn(15 downto 11) is
					when "10000" => -- ��Ȩָ��
						if Lf = '0' then
							case Insn(3 downto 0) is
								when "0000" => -- MTUP
									Reg1(3) <= '0';
									Reg1(2 downto 0) <= Insn(10 downto 8);
									RegDst <= "1101";
									RegWr <= '1';
								when "0001" => -- MTKP
									Reg1(3) <= '0';
									Reg1(2 downto 0) <= Insn(10 downto 8);
									RegDst <= "1100";
									RegWr <= '1';
								when "0010" => -- MFUP
									Reg1 <= "1101";
									RegDst(3) <= '0';
									RegDst(2 downto 0) <= Insn(10 downto 8);
									RegWr <= '1';
								when "0011" => -- MFKP
									Reg1 <= "1100";
									RegDst(3) <= '0';
									RegDst(2 downto 0) <= Insn(10 downto 8);
									RegWr <= '1';
								when "0100" => -- SVUP
									Reg1 <= "1000";
									RegDst <= "1101";
									RegWr <= '1';
								when "0101" => -- LDKP
									Reg1 <= "1100";
									RegDst <= "1000";
									RegWr <= '1';
								when "0110" => -- EJR
									Reg2(3) <= '0';
									Reg2(2 downto 0) <= Insn(10 downto 8);
									Jcond <= "110"; -- Data2
									Degrade <= '1'; -- �������м�
								when others => -- �Ƿ�ָ��
									Inval <= '1';
							end case;
						else -- ��Ȩ�쳣
							Priv <= '1';
						end if;
					when "11111" => -- INT
						Int <= '1';
					when "01001" => -- ADDIU
						Reg1(3) <= '0';
						Reg1(2 downto 0) <= Insn(10 downto 8); -- Reg1 <= Rx
						RegDst(3) <= '0'; 							-- RegDst <= Rx
						RegDst(2 downto 0) <= Insn(10 downto 8);
						-- �����������ֽ��з�����չ Imm <= SignExtend(Insn(7 downto 0))
						case Insn(7) is
							when '1' => Imm(15 downto 8) <= "11111111";
							when others => Imm(15 downto 8) <= "00000000";
						end case;
						Imm(7 downto 0) <= Insn(7 downto 0);
						Op2Src <= '1'; -- Imm
						RegWr <= '1'; -- Yes
					when "01000" => -- ADDIU3
						Reg1(3) <= '0'; -- Reg1 <= Rx
						Reg1(2 downto 0) <= Insn(10 downto 8);
						RegDst(3) <= '0'; -- RegDst <= Ry
						RegDst(2 downto 0) <= Insn(7 downto 5);
						-- �����������з�����չ Imm <= SignExtend(Insn(3 downto 0))
						case Insn(3) is
							when '1' => Imm(15 downto 4) <= "111111111111";
							when others => Imm(15 downto 4) <= "000000000000";
						end case;
						Imm(3 downto 0) <= Insn(3 downto 0);
						Op2Src <= '1'; -- Imm
						RegWr <= '1'; -- Yes
					when "11100" => -- ADDU/SUBU
						case Insn(1 downto 0) is
						 when "01" => -- ADDU
							Reg1(3) <= '0'; -- Reg1 <= Rx
							Reg1(2 downto 0) <= Insn(10 downto 8);
							Reg2(3) <= '0'; -- Reg2 <= Ry
							Reg2(2 downto 0) <= Insn(7 downto 5);
							RegDst(3) <= '0'; -- RegDst <= Rz
							RegDst(2 downto 0) <= Insn(4 downto 2);
							RegWr <= '1'; -- Yes
						 when "11" => -- SUBU
							Reg1(3) <= '0'; -- Reg1 <= Rx
							Reg1(2 downto 0) <= Insn(10 downto 8);
							Reg2(3) <= '0'; -- Reg2 <= Ry
							Reg2(2 downto 0) <= Insn(7 downto 5);
							RegDst(3) <= '0'; -- RegDst <= Rz
							RegDst(2 downto 0) <= Insn(4 downto 2);
							AluOp <= "0001"; -- Subtract
							RegWr <= '1'; -- Yes
						 when others => -- �Ƿ�ָ��
							Inval <= '1';
						end case;
					when "11101" => -- AND/JALR/JR/JRRA/MFPC/NEG/NOT/OR/CMP
						case Insn(4 downto 0) is
							when "01100" => -- AND
								Reg1(3) <= '0'; -- Reg1 <= Rx
								Reg1(2 downto 0) <= Insn(10 downto 8);
								Reg2(3) <= '0'; -- Reg2 <= Ry
								Reg2(2 downto 0) <= Insn(7 downto 5);
								RegDst(3) <= '0'; -- RegDst <= Rx
								RegDst(2 downto 0) <= Insn(10 downto 8);
								AluOp <= "0010"; -- AND(2)
								RegWr <= '1'; -- Yes
							when "01011" => -- NEG
								Reg2(3) <= '0'; -- Reg2 <= Ry
								Reg2(2 downto 0) <= Insn(7 downto 5);
								RegDst(3) <= '0'; -- RegDst <= Rx
								RegDst(2 downto 0) <= Insn(10 downto 8);
								AluOp <= "0101"; -- NEG
								RegWr <= '1'; -- Yes
							when "01111" => -- NOT
								Reg2(3) <= '0'; -- Reg2 <= Ry
								Reg2(2 downto 0) <= Insn(7 downto 5);
								RegDst(3) <= '0'; -- RegDst <= Rx
								RegDst(2 downto 0) <= Insn(10 downto 8);
								AluOp <= "0110"; -- NOT
								RegWr <= '1'; -- Yes
							when "01101" => -- OR
								Reg1(3) <= '0'; -- Reg1 <= Rx
								Reg1(2 downto 0) <= Insn(10 downto 8);
								Reg2(3) <= '0'; -- Reg2 <= Ry
								Reg2(2 downto 0) <= Insn(7 downto 5);
								RegDst(3) <= '0'; -- RegDst <= Rx
								RegDst(2 downto 0) <= Insn(10 downto 8);
								AluOp <= "0011"; -- Or
								RegWr <= '1'; -- Yes
							when "01010" => -- CMP
								Reg1(3) <= '0'; -- Reg1 <= Rx
								Reg1(2 downto 0) <= Insn(10 downto 8);
								Reg2(3) <= '0'; -- Reg2 <= Rx
								Reg2(2 downto 0) <= Insn(7 downto 5);
								RegDst <= "1111"; -- RegDst <= ZERO
								AluOp <= "0100"; -- (4) Equal test
								TWr <= '1'; -- Yes
							when "00000" => -- JALR/JR/JRRA/MFPC
								case Insn(7 downto 5) is
									when "110" => -- JALR
										Reg2(3) <= '0'; -- Reg2 <= Rx
										Reg2(2 downto 0) <= Insn(10 downto 8);
										RegDst <= "1010"; -- RegDst <= RA
										Op1Src <= '1'; -- PC
										Op2Src <= '1'; -- Imm
										Jcond <= "110"; -- ��������ת��PCֵ����Data2
										RegWr <= '1'; -- Yes
									when "000" => -- JR
										Reg2(3) <= '0'; -- Reg2 <= Rx
										Reg2(2 downto 0) <= Insn(10 downto 8);
										Jcond <= "110"; -- ��������ת��PCֵ����Data2
									when "001" => -- JRRA
										Reg2 <= "1010"; -- Reg2 <= RA
										Jcond <= "110"; -- ��������ת��PCֵ����Data2
									when "010" => -- MFPC
										RegDst(3) <= '0'; -- RegDst <= Rx
										RegDst(2 downto 0) <= Insn(10 downto 8);
										Op1Src <= '1'; -- PC
										RegWr <= '1'; -- Yes
									when others => -- �Ƿ�ָ��
										Inval <= '1';
								end case;
							when others => -- ����ָ��
								Inval <= '1';
						end case;
					when "00010" => -- B
						-- Imm <= SignExtend(Insn(10 downto 0))
						case Insn(10) is
							when '1' => Imm(15 downto 11) <= "11111";
							when others => Imm(15 downto 11) <= "00000";
						end case;
						Imm(10 downto 0) <= Insn(10 downto 0);
						Op1Src <= '1'; -- PC
						Op2Src <= '1'; -- Imm
						Jcond <= "001"; -- Unconditional jump
					when "00100" => -- BEQZ
						Reg2(3) <= '0'; -- Reg2 <= Rx
						Reg2(2 downto 0) <= Insn(10 downto 8);
						RegDst <= "1111"; -- RegDst <= ZERO
						-- Imm <= SignExtend(Insn(7 downto 0));
						case Insn(7) is
							when '1' => Imm(15 downto 8) <= "11111111";
							when others => Imm(15 downto 8) <= "00000000";
						end case;
						Imm(7 downto 0) <= Insn(7 downto 0);
						Op1Src <= '1'; -- PC
						Op2Src <= '1'; -- Imm
						Jcond <= "101"; -- (5) Jump if Data2 is zero (ZCMP == 1)
					when "00101" => -- BNEZ
						Reg2(3) <= '0'; -- Reg2 <= Rx
						Reg2(2 downto 0) <= Insn(10 downto 8);
						-- Imm <= SignExtend(Insn(7 downto 0));
						case Insn(7) is
							when '1' => Imm(15 downto 8) <= "11111111";
							when others => Imm(15 downto 8) <= "00000000";
						end case;
						Imm(7 downto 0) <= Insn(7 downto 0);
						Op1Src <= '1'; -- PC
						Op2Src <= '1'; -- Imm
						Jcond <= "100"; -- (4) Jump if Data2 is nonzero (ZCMP == 0)
					when "01100" => -- BTEQZ/BTNEZ/MTSP
						case Insn(10 downto 8) is
							when "011" => -- ADDSP
								Reg1 <= "1000"; -- Reg1 <= SP
								RegDst <= "1000"; -- RegDst <= SP
								-- Imm <= SignExtend(Insn(7 downto 0))
								case Insn(7) is
									when '1' => Imm(15 downto 8) <= "11111111";
									when others => Imm(15 downto 8) <= "00000000";
								end case;
								Imm(7 downto 0) <= Insn(7 downto 0);
								Op2Src <= '1'; -- Imm
								RegWr <= '1'; -- Yes
							when "000" => -- BTEQZ
								-- Imm <= SignExtend(Insn(7 downto 0))
								case Insn(7) is
									when '1' => Imm(15 downto 8) <= "11111111";
									when others => Imm(15 downto 8) <= "00000000";
								end case;
								Imm(7 downto 0) <= Insn(7 downto 0);
								Op1Src <= '1'; -- PC
								Op2Src <= '1'; -- Imm
								Jcond <= "010"; -- (2) Jump if T == 0
							when "001" => -- BTNEZ
								-- Imm <= SignExtend(Insn(7 downto 0))
								case Insn(7) is
									when '1' => Imm(15 downto 8) <= "11111111";
									when others => Imm(15 downto 8) <= "00000000";
								end case;
								Imm(7 downto 0) <= Insn(7 downto 0);
								Op1Src <= '1'; -- PC
								Op2Src <= '1'; -- Imm
								Jcond <= "011"; -- (3) Jump if T != 0
							when "100" => -- MTSP
								Reg1(3) <= '0'; -- Reg1 <= Ry
								Reg1(2 downto 0) <= Insn(7 downto 5);
								RegDst <= "1000"; -- RegDst <= SP
								RegWr <= '1'; -- Yes
							when others => -- �Ƿ�ָ��
								Inval <= '1';
						end case;
					when "01101" => -- LI
						RegDst(3) <= '0'; -- RegDst <= Rx
						RegDst(2 downto 0) <= Insn(10 downto 8);
						-- Imm <= ZeroExtend(Insn(7 downto 0))
						Imm(15 downto 8) <= "00000000";
						Imm(7 downto 0) <= Insn(7 downto 0);
						Op2Src <= '1'; -- Imm
						RegWr <= '1'; -- Yes
					when "10011" => -- LW
						Reg1(3) <= '0'; -- Reg1 <= Rx
						Reg1(2 downto 0) <= Insn(10 downto 8);
						RegDst(3) <= '0'; -- RegDst <= Ry
						RegDst(2 downto 0) <= Insn(7 downto 5);
						-- Imm <= SignExtend(Insn(4 downto 0))
						case Insn(4) is
							when '1' => Imm(15 downto 5) <= "11111111111";
							when others => Imm(15 downto 5) <= "00000000000";
						end case;
						Imm(4 downto 0) <= Insn(4 downto 0);
						Op2Src <= '1'; -- Imm
						MemRd <= '1'; -- Yes
						RegWr <= '1'; -- Yes
					when "10010" => -- LW_SP
						Reg1 <= "1000"; -- Reg1 <= SP
						RegDst(3) <= '0'; -- RegDst <= Rx
						RegDst(2 downto 0) <= Insn(10 downto 8);
						-- Imm <= SignExtend(Insn(7 downto 0))
						case Insn(7) is
							when '1' => Imm(15 downto 8) <= "11111111";
							when others => Imm(15 downto 8) <= "00000000";
						end case;
						Imm(7 downto 0) <= Insn(7 downto 0);
						Op2Src <= '1'; -- Imm
						MemRd <= '1'; -- Yes
						RegWr <= '1'; -- Yes
					when "11110" => -- MFIH/MTIH
						case Insn(7 downto 0) is
							when "00000000" => -- MFIH
								Reg1 <= "1001"; -- Reg1 <= IH
								RegDst(3) <= '0'; -- RegDst <= Rx
								RegDst(2 downto 0) <= Insn(10 downto 8);
								RegWr <= '1'; -- Yes
							when "00000001" => -- MTIH
								Reg1(3) <= '0'; -- Reg1 <= Rx
								Reg1(2 downto 0) <= Insn(10 downto 8);
								RegDst <= "1001"; -- RegDst <= IH
								RegWr <= '1'; -- Yes
							when others => -- �Ƿ�ָ��
								Inval <= '1';
						end case;
					when "00001" => -- NOP
					when "00110" => -- SLL/SRA
						case Insn(1 downto 0) is
							when "00" => -- SSL
								Reg1(3) <= '0'; -- Reg1 <= Ry
								Reg1(2 downto 0) <= Insn(7 downto 5);
								RegDst(3) <= '0'; -- RegDst <= Rx
								RegDst(2 downto 0) <= Insn(10 downto 8);
								-- Imm <= ZeroExtend(Insn(4 downto 2))
								Imm(15 downto 3) <= "0000000000000";
								Imm(2 downto 0) <= Insn(4 downto 2);
								Op2Src <= '1'; -- Imm
								AluOp <= "0111"; -- SLL
								RegWr <= '1'; -- Yes
							when "11" => -- SRA
								Reg1(3) <= '0'; -- Reg1 <= Ry
								Reg1(2 downto 0) <= Insn(7 downto 5);
								RegDst(3) <= '0'; -- RegDst <= Rx
								RegDst(2 downto 0) <= Insn(10 downto 8);
								-- Imm <= ZeroExtend(Insn(4 downto 2))
								Imm(15 downto 3) <= "0000000000000";
								Imm(2 downto 0) <= Insn(4 downto 2);
								Op2Src <= '1'; -- Imm
								AluOp <= "1000"; -- SLL
								RegWr <= '1'; -- Yes
							when others => --����ָ��
								Inval <= '1';
						end case;
					when "11011" => -- SW
						Reg1(3) <= '0'; -- Reg1 <= Rx
						Reg1(2 downto 0) <= Insn(10 downto 8);
						Reg2(3) <= '0'; -- Reg2 <= Ry
						Reg2(2 downto 0) <= Insn(7 downto 5);
						-- Imm <= SignExtend(Insn(4 downto 0))
						case Insn(4) is
							when '1' => Imm(15 downto 5) <= "11111111111";
							when others => Imm(15 downto 5) <= "00000000000";
						end case;
						Imm(4 downto 0) <= Insn(4 downto 0);
						Op2Src <= '1'; -- Imm
						MemWr <= '1'; -- Yes
					when "11010" => -- SW_SP
						Reg1 <= "1000"; -- Reg1 <= SP
						Reg2(3) <= '0'; -- Reg2 <= Rx
						Reg2(2 downto 0) <= Insn(10 downto 8);
						-- Imm <= SignExtend(Insn(7 downto 0))
						case Insn(7) is
							when '1' => Imm(15 downto 8) <= "11111111";
							when others => Imm(15 downto 8) <= "00000000";
						end case;
						Imm(7 downto 0) <= Insn(7 downto 0);
						Op2Src <= '1'; -- Imm
						MemWr <= '1'; -- Yes
					when others => -- �Ƿ�ָ��
						Inval <= '1';
				end case;
		end case;
	end process;
end Behavioral;

